module top ();
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C31 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C28 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_1uF_10V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C27 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C26 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C30 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C29 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_243R_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R7 ( .PIN1(GND), .PIN2(Net__R7_Pad2_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C22 ( .PIN2(S0SVREF), .PIN1(GND) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R3 ( .PIN1(S0SCK_P), .PIN2(Net__R3_Pad2_) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R4 ( .PIN1(S0SCK_N), .PIN2(Net__R4_Pad2_) );
  CELL_243R_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R9 ( .PIN2(GND), .PIN1(Net__R9_Pad1_) );
  NA_243R_1___OLIMEX_RLC_FP_R_0402_5MIL_DWS R13 ( .PIN2(GND), .PIN1(Net__R13_Pad1_) );
  CELL_2k_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R8 ( .PIN2(VREF0_DDR3), .PIN1(GND) );
  CELL_2k_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R5 ( .PIN2(_1_5V), .PIN1(VREF0_DDR3) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C11 ( .PIN1(_1_5V), .PIN2(VREF0_DDR3) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C23 ( .PIN1(VREF0_DDR3), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C24 ( .PIN1(VREF0_DDR3), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C12 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C13 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C14 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C15 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C16 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C1 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C2 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C3 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C4 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C5 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_2k_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R12 ( .PIN2(S0SVREF), .PIN1(GND) );
  CELL_2k_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R11 ( .PIN2(_1_5V), .PIN1(S0SVREF) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C32 ( .PIN2(_1_5V), .PIN1(S0SVREF) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C33 ( .PIN2(S0SVREF), .PIN1(GND) );
  CELL_243R_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R10 ( .PIN1(Net__R10_Pad1_), .PIN2(GND) );
  NA_243R_1___OLIMEX_RLC_FP_R_0402_5MIL_DWS R14 ( .PIN1(Net__R14_Pad1_), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C25 ( .PIN1(VREF0_DDR3), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C17 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C18 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C19 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C20 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C21 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C6 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C7 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C8 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C9 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C10 ( .PIN1(_1_5V), .PIN2(GND) );
  CELL_100R_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R2 ( .PIN1(S0SCK_N), .PIN2(S0SCK_P) );
  CELL_2k_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R1 ( .PIN2(_1_5V), .PIN1(S0SRST) );
  NA_OLIMEX_RLC_FP_R_0402_5MIL_DWS R6 ( .PIN2(S0SVREF), .PIN1(VREF0_DDR3) );
  K4B4G1646Q_HYK0_FBGA_96_256Mx16_DDR3_1600_11_11_11__OLIMEX_IC_FP_FBGA96_HYNIX_SAMSUNG_512MX16_DDR3_ U2 ( .N9(_1_5V), .R1(_1_5V), .R9(_1_5V), .A1(_1_5V), .A8(_1_5V), .B2(_1_5V), .G7(_1_5V), .C1(_1_5V), .H2(_1_5V), .H9(_1_5V), .C9(_1_5V), .D2(_1_5V), .D9(_1_5V), .E9(_1_5V), .F1(_1_5V), .K2(_1_5V), .K8(_1_5V), .N1(_1_5V), .T2(S0SRST), .K7(S0SCK_N), .J7(S0SCK_P), .M8(VREF0_DDR3), .H1(VREF0_DDR3), .D8(GND), .G9(GND), .B1(GND), .B3(GND), .B9(GND), .F9(GND), .G1(GND), .G8(GND), .A9(GND), .J2(GND), .D1(GND), .E1(GND), .E2(GND), .E8(GND), .P1(GND), .P9(GND), .T1(GND), .M1(GND), .M9(GND), .T9(GND), .J8(GND), .R2(S0SA7), .M2(S0SBA0), .M7(S0SA15), .T7(S0SA14), .T3(S0SA13), .N7(S0SA12), .R7(S0SA11), .L7(S0SA10), .R3(S0SA9), .T8(S0SA8), .R8(S0SA6), .P2(S0SA5), .P8(S0SA4), .N2(S0SA3), .P3(S0SA2), .P7(S0SA1), .N3(S0SA0), .L9(Net__R13_Pad1_), .L8(Net__R9_Pad1_), .A2(S0SDQ15), .C3(S0SDQ14), .C2(S0SDQ13), .A3(S0SDQ12), .N8(S0SBA1), .J1(S0SODT1), .K1(S0SODT0), .J3(S0SRAS), .K3(S0SCAS), .L3(S0SWE), .L1(S0SCS1), .L2(S0SCS0), .J9(S0SCKE1), .K9(S0SCKE0), .M3(S0SBA2), .D7(S0SDQ11), .B8(S0SDQ10), .C8(S0SDQ9), .A7(S0SDQ8), .F8(S0SDQ7), .H8(S0SDQ6), .H3(S0SDQ5), .E3(S0SDQ4), .H7(S0SDQ3), .F2(S0SDQ2), .G2(S0SDQ1), .F7(S0SDQ0), .F3(S0SDQS0_P), .B7(S0SDQS1_N), .C7(S0SDQS1_P), .D3(S0SDQM1), .E7(S0SDQM0), .G3(S0SDQS0_N) );
  K4B4G1646Q_HYK0_FBGA_96_256Mx16_DDR3_1600_11_11_11__OLIMEX_IC_FP_FBGA96_HYNIX_SAMSUNG_512MX16_DDR3_ U3 ( .N9(_1_5V), .R1(_1_5V), .R9(_1_5V), .K8(_1_5V), .N1(_1_5V), .G7(_1_5V), .H2(_1_5V), .H9(_1_5V), .K2(_1_5V), .A8(_1_5V), .B2(_1_5V), .C1(_1_5V), .A1(_1_5V), .C9(_1_5V), .D2(_1_5V), .D9(_1_5V), .E9(_1_5V), .F1(_1_5V), .T2(S0SRST), .K7(S0SCK_N), .J7(S0SCK_P), .H1(VREF0_DDR3), .M8(VREF0_DDR3), .L9(Net__R14_Pad1_), .L8(Net__R10_Pad1_), .M9(GND), .M1(GND), .G8(GND), .D8(GND), .D1(GND), .E1(GND), .E2(GND), .E8(GND), .F9(GND), .A9(GND), .B3(GND), .B9(GND), .B1(GND), .G9(GND), .J2(GND), .J8(GND), .P1(GND), .P9(GND), .T1(GND), .T9(GND), .G1(GND), .R2(S0SA7), .M2(S0SBA0), .M7(S0SA15), .T7(S0SA14), .T3(S0SA13), .N7(S0SA12), .R7(S0SA11), .L7(S0SA10), .R3(S0SA9), .T8(S0SA8), .R8(S0SA6), .P2(S0SA5), .P8(S0SA4), .N2(S0SA3), .P3(S0SA2), .P7(S0SA1), .N3(S0SA0), .N8(S0SBA1), .F8(S0SDQ19), .H7(S0SDQ18), .H8(S0SDQ17), .F7(S0SDQ16), .H3(S0SDQ20), .A2(S0SDQ30), .C2(S0SDQ31), .C3(S0SDQ29), .A3(S0SDQ28), .B8(S0SDQ27), .D7(S0SDQ26), .C8(S0SDQ25), .A7(S0SDQ24), .G2(S0SDQ23), .E3(S0SDQ22), .F2(S0SDQ21), .F3(S0SDQS2_P), .J1(S0SODT1), .K1(S0SODT0), .J3(S0SRAS), .K3(S0SCAS), .L3(S0SWE), .L1(S0SCS1), .L2(S0SCS0), .G3(S0SDQS2_N), .B7(S0SDQS3_N), .C7(S0SDQS3_P), .D3(S0SDQM3), .E7(S0SDQM2), .J9(S0SCKE1), .K9(S0SCKE0), .M3(S0SBA2) );
  AllWinner_A64_FBGA396__OLIMEX_IC_FP_FBGA396 U1 ( .G7(_1_5V), .G8(_1_5V), .J8(_1_5V), .G9(_1_5V), .K6(_1_5V), .K7(_1_5V), .L6(_1_5V), .N8(_1_5V), .L8(_1_5V), .N7(_1_5V), .L7(_1_5V), .D10(S0SRST), .G5(S0SVREF), .J15(GND), .P11(GND), .P12(GND), .P13(GND), .V8(GND), .M8(GND), .M9(GND), .N10(GND), .N11(GND), .N12(GND), .N13(GND), .P7(GND), .N15(GND), .N4(GND), .N9(GND), .P10(GND), .U11(GND), .U12(GND), .T13(GND), .M3(GND), .T8(GND), .T9(GND), .R5(GND), .P9(GND), .R10(GND), .R11(GND), .R12(GND), .R6(GND), .R7(GND), .R8(GND), .R9(GND), .T10(GND), .T11(GND), .T12(GND), .R15(GND), .P8(GND), .V14(GND), .U2(GND), .U5(GND), .U7(GND), .U8(GND), .U9(GND), .K8(GND), .K9(GND), .L10(GND), .L11(GND), .AC23(GND), .A1(GND), .C3(GND), .C7(GND), .A23(GND), .L12(GND), .M15(GND), .K12(GND), .J14(GND), .J9(GND), .K10(GND), .K11(GND), .J11(GND), .K13(GND), .D7(GND), .L4(GND), .L5(GND), .L9(GND), .M10(GND), .M11(GND), .M12(GND), .L15(GND), .G11(GND), .G6(GND), .H13(GND), .H4(GND), .J10(GND), .E4(S0SA7), .D8(S0SBA0), .T4(S0SA15), .K4(S0SA14), .E8(S0SA13), .K5(S0SA12), .U4(S0SA11), .M4(S0SA10), .C4(S0SA9), .D3(S0SA8), .F3(S0SA6), .G4(S0SA5), .P6(S0SA4), .N6(S0SA3), .N5(S0SA2), .R4(S0SA1), .P5(S0SA0), .M2(S0SDQ15), .N1(S0SDQ14), .N2(S0SDQ13), .N3(S0SDQ12), .R3(S0SBA1), .E1(S0SDQ19), .E2(S0SDQ18), .F2(S0SDQ17), .E3(S0SDQ16), .B1(S0SDQ20), .B8(S0SDQ30), .B9(S0SDQ31), .A8(S0SDQ29), .A7(S0SDQ28), .A5(S0SDQ27), .A4(S0SDQ26), .B4(S0SDQ25), .C5(S0SDQ24), .B3(S0SDQ23), .A2(S0SDQ22), .B2(S0SDQ21), .D2(S0SDQS2_P), .E7(S0SODT1), .D5(S0SODT0), .F7(S0SRAS), .C9(S0SCAS), .C8(S0SWE), .H5(S0SCS1), .E5(S0SCS0), .D1(S0SDQS2_N), .B5(S0SDQS3_N), .B6(S0SDQS3_P), .B7(S0SDQM3), .C2(S0SDQM2), .H6(S0SCKE1), .J3(S0SCKE0), .C6(S0SBA2), .R2(S0SDQ11), .T1(S0SDQ10), .T2(S0SDQ9), .T3(S0SDQ8), .L2(S0SDQ7), .L1(S0SDQ6), .H1(S0SDQ5), .H2(S0SDQ4), .K1(S0SDQ3), .H3(S0SDQ2), .U1(Net__R7_Pad2_), .G1(S0SDQ1), .L3(S0SDQ0), .K3(S0SDQS0_P), .P2(S0SDQS1_N), .P1(S0SDQS1_P), .P3(S0SDQM1), .J2(S0SDQM0), .K2(S0SDQS0_N), .G3(Net__R4_Pad2_), .G2(Net__R3_Pad2_), .N19(_3_3V), .L16(_3_3V), .T14(_3_3V), .U15(_3_3V), .U16(_3_3V), .N18(_3_3V), .G13(Net__C54_Pad2_), .F12(Net__C54_Pad2_), .E11(Net__C61_Pad1_), .E10(Net__C61_Pad2_), .E13(_1_8V), .B11(Net__C59_Pad1_), .B12(Net__C55_Pad1_), .C11(Net__C51_Pad1_), .N16(_3_0VA), .G14(_3_0VA), .A11(GNDA), .D13(Net__C63_Pad1_), .K18(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_ALE_SDC2_DS), .T21(SPI0_MOSI), .R16(VCC_PC), .E14(NAND_Flash___eMMC__T_Card_and_Audio_MBIAS), .B15(NAND_Flash___eMMC__T_Card_and_Audio_MICIN1P), .B17(NAND_Flash___eMMC__T_Card_and_Audio_MICIN2P), .E16(Net__U1_PadE16_), .F16(Net__U1_PadF16_), .C14(Net__U1_PadC14_), .D14(Net__U1_PadD14_), .B13(Net__U1_PadB13_), .A13(Net__U1_PadA13_), .B10(Net__U1_PadB10_), .C12(NAND_Flash___eMMC__T_Card_and_Audio_HPOUTR), .C10(NAND_Flash___eMMC__T_Card_and_Audio_HPOUTFB), .B16(NAND_Flash___eMMC__T_Card_and_Audio_MICIN1N), .D11(NAND_Flash___eMMC__T_Card_and_Audio_HP_DET), .M21(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ0_SDC2_D0), .L19(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ1_SDC2_D1), .K20(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ2_SDC2_D2), .H20(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ3_SDC2_D3), .P18(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ4_SDC2_D4), .L20(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ5_SDC2_D5), .J21(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ6_SDC2_D6), .R21(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ7_SDC2_D7), .N20(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQS_SDC2_RST), .G20(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_RE_SDC2_CLK), .K19(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_RB0_SDC2_CMD), .P20(SPI0_CLK), .P19(SPI0_CS), .T20(PC4), .T19(PC7), .AB9(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D2), .AC8(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_CLK), .W9(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_CMD), .AB8(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_DET_), .AB6(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D3), .AB10(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D1), .W13(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D0), .C16(NAND_Flash___eMMC__T_Card_and_Audio_LINEOUTR), .D16(NAND_Flash___eMMC__T_Card_and_Audio_LINEOUTL), .C13(NAND_Flash___eMMC__T_Card_and_Audio_HPOUTL), .A17(NAND_Flash___eMMC__T_Card_and_Audio_MICIN2N), .A14(NAND_Flash___eMMC__T_Card_and_Audio_LINEINR), .B14(NAND_Flash___eMMC__T_Card_and_Audio_LINEINL), .H16(net_3_0V_RTC), .H19(Net__HSIC1_Pad2_), .G19(Net__HSIC1_Pad3_), .T23(Power_Supply__Extensions_and_MiPi_DSI_DSI_D0N), .D22(PL12), .C19(PL7), .B21(PL8), .D20(PL9), .D21(PL10), .C20(PL11), .F17(UBOOT), .Y22(Power_Supply__Extensions_and_MiPi_DSI_PE13), .AA21(Power_Supply__Extensions_and_MiPi_DSI_PE3), .AA22(Power_Supply__Extensions_and_MiPi_DSI_PE2), .AB23(Power_Supply__Extensions_and_MiPi_DSI_PE1), .AA18(Power_Supply__Extensions_and_MiPi_DSI_PE0), .W22(Power_Supply__Extensions_and_MiPi_DSI_PE17_GPIO_LED), .AB21(Power_Supply__Extensions_and_MiPi_DSI_PE16), .Y23(Power_Supply__Extensions_and_MiPi_DSI_PE15), .AC20(Power_Supply__Extensions_and_MiPi_DSI_PE14), .AA19(Power_Supply__Extensions_and_MiPi_DSI_PE4), .AB20(Power_Supply__Extensions_and_MiPi_DSI_PE12), .W21(Power_Supply__Extensions_and_MiPi_DSI_PE11), .AB22(Power_Supply__Extensions_and_MiPi_DSI_PE10), .Y17(Power_Supply__Extensions_and_MiPi_DSI_PE9), .AC22(Power_Supply__Extensions_and_MiPi_DSI_PE8), .Y19(Power_Supply__Extensions_and_MiPi_DSI_PE7), .W20(Power_Supply__Extensions_and_MiPi_DSI_PE6), .W17(Power_Supply__Extensions_and_MiPi_DSI_PE5), .AA7(Power_Supply__Extensions_and_MiPi_DSI_PB3), .W10(Power_Supply__Extensions_and_MiPi_DSI_PB2), .AB7(Power_Supply__Extensions_and_MiPi_DSI_PB1), .V9(Power_Supply__Extensions_and_MiPi_DSI_PB0), .AA6(Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_RST), .W8(Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_BKL), .Y6(Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_EN), .L22(Power_Supply__Extensions_and_MiPi_DSI_DSI_D3N), .E17(AP_RESET_), .W7(Power_Supply__Extensions_and_MiPi_DSI_PB4), .U18(Net__3_3V_VCC_PE_2_8V1_Pad2_), .A16(KEYADC), .P16(Net__C188_Pad2_), .H14(Net__R96_Pad1_), .AA11(Net__R97_Pad1_), .AA12(Net__R98_Pad1_), .G16(Net__C192_Pad2_), .V10(Net__DBG_UART1_Pad1_), .T17(_3_3VWiFiIO), .B18(AP_CK32KO), .K22(Net__C187_Pad1_), .K23(Net__R94_Pad1_), .B19(Net__C183_Pad1_), .C18(Net__C184_Pad1_), .W11(TWI0_SCK), .AB5(UART3_TX), .H15(net_1_1V_CPUS), .C17(PMU_SDA), .J16(VCC_PL), .T6(VDDFB_CPUX), .AC7(UART3_RX), .AA9(TWI1_SDA), .N23(Power_Supply__Extensions_and_MiPi_DSI_DSI_CKP), .L23(Power_Supply__Extensions_and_MiPi_DSI_DSI_D3P), .N22(Power_Supply__Extensions_and_MiPi_DSI_DSI_D2N), .M22(Power_Supply__Extensions_and_MiPi_DSI_DSI_D2P), .R22(Power_Supply__Extensions_and_MiPi_DSI_DSI_D1N), .P22(Power_Supply__Extensions_and_MiPi_DSI_DSI_D1P), .T22(Power_Supply__Extensions_and_MiPi_DSI_DSI_D0P), .P23(Power_Supply__Extensions_and_MiPi_DSI_DSI_CKN), .AA10(TWI0_SDA), .K16(net_1_2V_HSIC), .M16(_3_3VD), .AC4(TWI1_SCK), .Y7(Net__D4_Pad2_), .T15(net_1_1V_SYS), .J12(net_1_1V_SYS), .J13(net_1_1V_SYS), .K14(net_1_1V_SYS), .M14(net_1_1V_SYS), .M13(net_1_1V_SYS), .L14(net_1_1V_SYS), .L13(net_1_1V_SYS), .N14(net_1_1V_SYS), .P14(net_1_1V_SYS), .R14(net_1_1V_SYS), .R13(net_1_1V_SYS), .AB2(net_1_1V_CPUX), .AA3(net_1_1V_CPUX), .AA1(net_1_1V_CPUX), .AC1(net_1_1V_CPUX), .AC2(net_1_1V_CPUX), .U6(net_1_1V_CPUX), .Y4(net_1_1V_CPUX), .Y3(net_1_1V_CPUX), .W5(net_1_1V_CPUX), .W4(net_1_1V_CPUX), .W3(net_1_1V_CPUX), .W1(net_1_1V_CPUX), .V6(net_1_1V_CPUX), .V5(net_1_1V_CPUX), .Y2(net_1_1V_CPUX), .V4(net_1_1V_CPUX), .V2(net_1_1V_CPUX), .V3(net_1_1V_CPUX), .Y8(PH10), .D17(PMU_SCK), .G18(AP_NMI_), .U21(USB1_DRV), .Y14(USB_HDMI_WiFi_BT_Ethernet_LCD_EPHY_RST_), .Y16(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD0_LCD_D15), .W16(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD1_LCD_D14), .AA13(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD2_LCD_D13), .V17(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD3_LCD_D12), .AB16(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCTL_LCD_D19), .Y13(USB_HDMI_WiFi_BT_Ethernet_LCD_GMDC_LCD_PWM), .AC10(USB_HDMI_WiFi_BT_Ethernet_LCD_GMDIO_LCD_PWR), .AB4(USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_VBUSDET), .A22(USB0_D_P), .B22(USB0_D_N), .AA8(USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_ID), .C22(USB_HDMI_WiFi_BT_Ethernet_LCD_USB1_DM), .B23(USB_HDMI_WiFi_BT_Ethernet_LCD_USB1_DP), .D23(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2P), .AB15(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D20), .Y11(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D10), .AA16(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D11), .AA20(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D2), .AA17(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D3), .W19(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D4), .AA14(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D5), .V18(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D6), .AA15(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D7), .A20(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_RST_N), .AB17(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_RX), .E21(USB_HDMI_WiFi_BT_Ethernet_LCD_HHPD), .AA5(PH11), .E20(USB_HDMI_WiFi_BT_Ethernet_LCD_HSDA), .E22(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2N), .E23(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1P), .F21(USB_HDMI_WiFi_BT_Ethernet_LCD_HCEC), .F22(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1N), .G21(USB_HDMI_WiFi_BT_Ethernet_LCD_HSCL), .G22(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0P), .G23(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0N), .H22(USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCP), .H23(USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCN), .AC5(USB_HDMI_WiFi_BT_Ethernet_LCD_PH7_CTP_INT), .Y10(USB_HDMI_WiFi_BT_Ethernet_LCD_PH8_CTP_RST), .B20(USB_HDMI_WiFi_BT_Ethernet_LCD_AP_WAKE_BT), .D19(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_WAKE_AP), .V21(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_CLK), .U20(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_CMD), .A19(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_PMU_EN), .E19(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_WAKE_AP), .U23(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_TX), .AC17(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_CTS), .AB19(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_SYNC), .AB18(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_CLK), .AC19(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_DIN), .U22(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_DOUT), .U19(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D0), .V22(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D1), .W23(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D3), .Y21(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D2), .AC11(USB_HDMI_WiFi_BT_Ethernet_LCD_GCLKIN_LCD_VSYNC), .AB12(Net__R19_Pad1_), .AC16(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCK_LCD_D18), .AB11(Net__R72_Pad1_), .AB14(Net__RM1_Pad4_2_), .AC13(Net__RM1_Pad1_2_), .AC14(Net__RM1_Pad3_2_), .AB13(Net__RM1_Pad2_2_) );
  NA_100nF_10V_10___OLIMEX_RLC_FP_C_0402_5MIL_DWS C37 ( .PIN1(GND), .PIN2(Net__C37_Pad2_) );
  NA_2_2uF_6_3V_10___OLIMEX_RLC_FP_C_0603_5MIL_DWS C38 ( .PIN1(GND), .PIN2(Net__C37_Pad2_) );
  NA_2_2uF_6_3V_10___OLIMEX_RLC_FP_C_0603_5MIL_DWS C36 ( .PIN1(GND), .PIN2(VCC_PC) );
  NA_100nF_10V_10___OLIMEX_RLC_FP_C_0402_5MIL_DWS C35 ( .PIN1(GND), .PIN2(VCC_PC) );
  NA_2_2uF_6_3V_10___OLIMEX_RLC_FP_C_0603_5MIL_DWS C43 ( .PIN2(GND), .PIN1(Net__C42_Pad1_) );
  NA_100nF_10V_10___OLIMEX_RLC_FP_C_0402_5MIL_DWS C44 ( .PIN2(GND), .PIN1(Net__C42_Pad1_) );
  NA_FB0805_600R_2A__OLIMEX_RLC_FP_L_0805_5MIL_DWS L1 ( .PIN1(_3_3V), .PIN2(Net__C42_Pad1_) );
  NA_22uF_6_3V_20___OLIMEX_RLC_FP_C_0603_5MIL_DWS C42 ( .PIN2(GND), .PIN1(Net__C42_Pad1_) );
  NA_10k__OLIMEX_RLC_FP_R_0402_5MIL_DWS R21 ( .PIN2(VCC_PC), .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_RB0_SDC2_CMD) );
  NA_10k__OLIMEX_RLC_FP_R_0402_5MIL_DWS R23 ( .PIN2(VCC_PC), .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQS_SDC2_RST) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C34 ( .PIN1(GND), .PIN2(VCC_PC) );
  MICRO_SD_TFC_WPAPR_08__OLIMEX_Connectors_FP_TFC_WPAPR_08 MICRO_SD1 ( .PIN10(GND), .PIN11(GND), .PIN6(GND), .PIN13(GND), .PIN12(GND), .PIN4(Net__C64_Pad1_), .PIN5(Net__MICRO_SD1_Pad5_), .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D2), .PIN3(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_CMD), .PIN9(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_DET_), .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D3), .PIN8(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D1), .PIN7(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D0) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R33 ( .PIN1(Net__MICRO_SD1_Pad5_), .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_CLK) );
  CELL_47uF_6_3V_20__OLIMEX_RLC_FP_C_0805_5MIL_DWS C64 ( .PIN2(GND), .PIN1(Net__C64_Pad1_) );
  FB0805_600R_2A_OLIMEX_RLC_FP_L_0805_5MIL_DWS L2 ( .PIN2(Net__C64_Pad1_), .PIN1(_3_3V) );
  RA1206__4x0603__4B8_100k_OLIMEX_RLC_FP_RA1206__4X0603__4B8_xx RM7 ( .PIN3_1(_3_3V), .PIN2_1(_3_3V), .PIN4_1(_3_3V), .PIN1_1(_3_3V), .PIN4_2(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D2), .PIN3_2(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_DET_), .PIN2_2(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D1), .PIN1_2(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D0) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R31 ( .PIN2(_3_3V), .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_CMD) );
  CELL_100k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R30 ( .PIN2(_3_3V), .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_SDC0_D3) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C46 ( .PIN1(_3_0VA), .PIN2(GNDA) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C49 ( .PIN1(_3_0VA), .PIN2(GNDA) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C51 ( .PIN1(Net__C51_Pad1_), .PIN2(GNDA) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C53 ( .PIN1(Net__C51_Pad1_), .PIN2(GNDA) );
  CELL_1uF_10V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C55 ( .PIN1(Net__C55_Pad1_), .PIN2(GNDA) );
  CELL_200k_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R27 ( .PIN1(Net__C59_Pad1_), .PIN2(GNDA) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C59 ( .PIN1(Net__C59_Pad1_), .PIN2(GNDA) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C63 ( .PIN2(GNDA), .PIN1(Net__C63_Pad1_) );
  SCJ325P00XG0B02G_OLIMEX_Connectors_FP_SCJ325P00XG0B02G MIC_LINEIN1 ( .PIN3(Net__LINEINR_MICIN1_Pad2_), .PIN1(Net__LINEINL_MICIN2_Pad2_), .PIN2(GNDA), .PIN4(Net__MIC_LINEIN1_Pad4_), .PIN5(Net__MIC_LINEIN1_Pad5_) );
  CELL_33pF_50V_5__OLIMEX_RLC_FP_C_0402_5MIL_DWS C48 ( .PIN1(GNDA), .PIN2(Net__C48_Pad2_) );
  CELL_33pF_50V_5__OLIMEX_RLC_FP_C_0402_5MIL_DWS C62 ( .PIN2(GNDA), .PIN1(Net__C62_Pad1_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C52 ( .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_MICIN1P), .PIN1(Net__C52_Pad1_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C60 ( .PIN1(Net__C60_Pad1_), .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_MICIN2P) );
  CELL_2k_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R26 ( .PIN1(Net__C60_Pad1_), .PIN2(Net__C57_Pad2_) );
  CELL_470R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R25 ( .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_MBIAS), .PIN1(Net__C57_Pad2_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C57 ( .PIN1(GNDA), .PIN2(Net__C57_Pad2_) );
  CELL_2k_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R29 ( .PIN2(Net__C57_Pad2_), .PIN1(Net__C52_Pad1_) );
  SCJ325P00XG0B02G_OLIMEX_Connectors_FP_SCJ325P00XG0B02G HEADPHONES_LINEOUT1 ( .PIN4(Net__HEADPHONES_LINEOUT1_Pad4_), .PIN5(Net__HEADPHONES_LINEOUT1_Pad5_), .PIN3(Net__HEADPHONES_LINEOUT1_Pad3_), .PIN2(Net__HEADPHONES_LINEOUT1_Pad2_), .PIN1(Net__HEADPHONES_LINEOUT1_Pad1_) );
  FB0805_600R_2A_OLIMEX_RLC_FP_L_0805_5MIL_DWS L3 ( .PIN1(Net__HPHONEOUTR_LINEOUTR1_Pad2_), .PIN2(Net__HEADPHONES_LINEOUT1_Pad3_) );
  FB0805_600R_2A_OLIMEX_RLC_FP_L_0805_5MIL_DWS L4 ( .PIN2(Net__HEADPHONES_LINEOUT1_Pad2_), .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_HPOUTFB) );
  FB0805_600R_2A_OLIMEX_RLC_FP_L_0805_5MIL_DWS L5 ( .PIN2(Net__HEADPHONES_LINEOUT1_Pad1_), .PIN1(Net__HPHONEOUTL_LINEOUTL1_Pad2_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C65 ( .PIN1(GNDA), .PIN2(Net__C65_Pad2_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C66 ( .PIN1(GNDA), .PIN2(Net__C66_Pad2_) );
  CELL_100k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R35 ( .PIN1(GNDA), .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_HPOUTR) );
  NA_1M__OLIMEX_RLC_FP_R_0402_5MIL_DWS R32 ( .PIN1(Net__HEADPHONES_LINEOUT1_Pad4_), .PIN2(_3_0VA) );
  CELL_0R_Board_Mounted__OLIMEX_RLC_FP_R_0402_5MIL_0R_Board_Mounted_ R34 ( .PIN1(GNDA), .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_HPOUTFB) );
  CELL_2_2uF_6_3V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C61 ( .PIN1(Net__C61_Pad1_), .PIN2(Net__C61_Pad2_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C54 ( .PIN2(Net__C54_Pad2_), .PIN1(GNDA) );
  CELL_2_2uF_6_3V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C56 ( .PIN2(Net__C54_Pad2_), .PIN1(GNDA) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C50 ( .PIN2(_1_8V), .PIN1(GNDA) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C47 ( .PIN2(_1_8V), .PIN1(GNDA) );
  CELL_0R_Board_Mounted__OLIMEX_RLC_FP_R_0603_5MIL_0R_Board_Mounted_ R36 ( .PIN1(GND), .PIN2(GNDA) );
  NA_W25Q128FVSIG__OLIMEX_IC_FP_SO_8_208mil U12 ( .PIN4(GND), .PIN8(_3_3V), .PIN5(SPI0_MOSI), .PIN2(SPI0_MISO), .PIN3(Net__R55_Pad1_), .PIN6(SPI0_CLK), .PIN1(SPI0_CS), .PIN7(Net__R57_Pad1_) );
  NA_100nF_10V_10___OLIMEX_RLC_FP_C_0402_5MIL_DWS C81 ( .PIN1(GND), .PIN2(_3_3V) );
  NA_10k__OLIMEX_RLC_FP_R_0402_5MIL_DWS R57 ( .PIN2(_3_3V), .PIN1(Net__R57_Pad1_) );
  NA_10k__OLIMEX_RLC_FP_R_0402_5MIL_DWS R56 ( .PIN2(_3_3V), .PIN1(Net__R55_Pad1_) );
  NA_OLIMEX_RLC_FP_R_0402_5MIL_DWS R55 ( .PIN2(GND), .PIN1(Net__R55_Pad1_) );
  NA_10k__OLIMEX_RLC_FP_R_0402_5MIL_DWS R53 ( .PIN2(_3_3V), .PIN1(SPI0_CS) );
  Opened_2_3__Soldered_1_2__OLIMEX_Jumpers_FP_SJ_2_SMALL LINEINR_MICIN1 ( .PIN2(Net__LINEINR_MICIN1_Pad2_), .PIN3(Net__C45_Pad1_), .PIN1(Net__C52_Pad1_) );
  Opened_2_3__Soldered_1_2__OLIMEX_Jumpers_FP_SJ_2_SMALL LINEINL_MICIN2 ( .PIN2(Net__LINEINL_MICIN2_Pad2_), .PIN1(Net__C60_Pad1_), .PIN3(Net__C58_Pad1_) );
  CELL_47k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R59 ( .PIN1(Net__HEADPHONES_LINEOUT1_Pad4_), .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_HP_DET) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R63 ( .PIN1(Net__C65_Pad2_), .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_HPOUTL) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R64 ( .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_HPOUTR), .PIN1(Net__C66_Pad2_) );
  Soldered_1_2__Opened_2_3__OLIMEX_Jumpers_FP_SJ_2_SMALL HPHONEOUTR_LINEOUTR1 ( .PIN2(Net__HPHONEOUTR_LINEOUTR1_Pad2_), .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_HPOUTR), .PIN3(Net__C86_Pad2_) );
  Soldered_1_2__Opened_2_3__OLIMEX_Jumpers_FP_SJ_2_SMALL HPHONEOUTL_LINEOUTL1 ( .PIN3(Net__C87_Pad2_), .PIN2(Net__HPHONEOUTL_LINEOUTL1_Pad2_), .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_HPOUTL) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C45 ( .PIN1(Net__C45_Pad1_), .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_LINEINR) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C58 ( .PIN1(Net__C58_Pad1_), .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_LINEINL) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C82 ( .PIN1(Net__C48_Pad2_), .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_MICIN1N) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C83 ( .PIN1(Net__C62_Pad1_), .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_MICIN2N) );
  CELL_33pF_50V_5__OLIMEX_RLC_FP_C_0402_5MIL_DWS C84 ( .PIN2(Net__C48_Pad2_), .PIN1(Net__C52_Pad1_) );
  CELL_33pF_50V_5__OLIMEX_RLC_FP_C_0402_5MIL_DWS C85 ( .PIN1(Net__C60_Pad1_), .PIN2(Net__C62_Pad1_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C86 ( .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_LINEOUTR), .PIN2(Net__C86_Pad2_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C87 ( .PIN2(Net__C87_Pad2_), .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_LINEOUTL) );
  TESTPAD_OLIMEX_Other_FP_TESTPAD_40_ROUND GNDA1 ( .PIN1(GNDA) );
  Mounting_hole_OLIMEX_Other_FP_Mounting_hole_3_3mm_with_5_5mm_pad Mounting_hole1 ( .PIN0(GND) );
  Mounting_hole_OLIMEX_Other_FP_Mounting_hole_3_3mm_with_5_5mm_pad Mounting_hole2 ( .PIN0(GND) );
  Mounting_hole_OLIMEX_Other_FP_Mounting_hole_3_3mm_with_5_5mm_pad Mounting_hole3 ( .PIN0(GND) );
  NA_KLMAG2GEND_B031_FBGA153___OLIMEX_IC_FP_FBGA153_Pitch_0_5mm_Ball_0_25mm_Dimensions_11_50x13_00x0_80mm U5 ( .P4(GND), .P6(GND), .K8(GND), .N2(GND), .N5(GND), .E7(GND), .G5(GND), .H10(GND), .J5(GND), .C4(GND), .A6(GND), .C2(Net__C37_Pad2_), .H5(Net__R15_Pad1_), .M6(NAND_Flash___eMMC__T_Card_and_Audio_eMMC_CLK), .J10(Net__C42_Pad1_), .F5(Net__C42_Pad1_), .E6(Net__C42_Pad1_), .K9(Net__C42_Pad1_), .P5(VCC_PC), .P3(VCC_PC), .N4(VCC_PC), .M4(VCC_PC), .C6(VCC_PC), .A3(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ0_SDC2_D0), .A4(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ1_SDC2_D1), .A5(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ2_SDC2_D2), .B2(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ3_SDC2_D3), .B3(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ4_SDC2_D4), .B4(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ5_SDC2_D5), .B5(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ6_SDC2_D6), .B6(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ7_SDC2_D7), .K5(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQS_SDC2_RST), .M5(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_RB0_SDC2_CMD) );
  NA_10k__OLIMEX_RLC_FP_R_0402_5MIL_DWS R67 ( .PIN2(VCC_PC), .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_DQ0_SDC2_D0) );
  Opened_OLIMEX_Jumpers_FP_SJ WP_Enable1 ( .PIN1(GND), .PIN2(Net__R55_Pad1_) );
  NA_22R__OLIMEX_RLC_FP_R_0402_5MIL_DWS R68 ( .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_eMMC_CLK), .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_RE_SDC2_CLK) );
  NA_OLIMEX_RLC_FP_C_0402_5MIL_DWS C94 ( .PIN2(GND), .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_eMMC_CLK) );
  CELL_0R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R66 ( .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_ALE_SDC2_DS), .PIN1(SPI0_MISO) );
  NA_10k__OLIMEX_RLC_FP_R_0402_5MIL_DWS R62 ( .PIN2(GND), .PIN1(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_ALE_SDC2_DS) );
  NA_22R__OLIMEX_RLC_FP_R_0402_5MIL_DWS R15 ( .PIN1(Net__R15_Pad1_), .PIN2(NAND_Flash___eMMC__T_Card_and_Audio_NAND0_ALE_SDC2_DS) );
  HDMI_SWM_19_OLIMEX_Connectors_FP_HDMI_SWM_19_Paste HDMI1 ( .PIN0(GND), .PIN5(GND), .PIN0(GND), .PIN0(GND), .PIN0(GND), .PIN11(GND), .PIN17(GND), .PIN2(GND), .PIN8(GND), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2P), .PIN13(Net__FET1_Pad3_), .PIN14(Net__HDMI1_Pad14_), .PIN19(Net__HDMI1_Pad19_), .PIN16(USB_HDMI_WiFi_BT_Ethernet_LCD_HSDA), .PIN3(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2N), .PIN4(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1P), .PIN6(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1N), .PIN15(USB_HDMI_WiFi_BT_Ethernet_LCD_HSCL), .PIN7(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0P), .PIN9(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0N), .PIN10(USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCP), .PIN12(USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCN), .PIN18(Net__D3_Pad1_) );
  NA_RCLAMP0524P_SLP2510P8___OLIMEX_IC_FP_SLP2510P8_TEST U7 ( .PIN3(GND), .PIN8(GND), .PIN10(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2P), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2P), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2N), .PIN9(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2N), .PIN4(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1P), .PIN7(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1P), .PIN6(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1N), .PIN5(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1N) );
  NA_RCLAMP0524P_SLP2510P8___OLIMEX_IC_FP_SLP2510P8_TEST U8 ( .PIN3(GND), .PIN8(GND), .PIN10(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0P), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0P), .PIN9(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0N), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0N), .PIN4(USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCP), .PIN7(USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCP), .PIN5(USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCN), .PIN6(USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCN) );
  NA_RCLAMP0524P_SLP2510P8___OLIMEX_IC_FP_SLP2510P8_TEST U10 ( .PIN3(GND), .PIN8(GND), .PIN6(USB_HDMI_WiFi_BT_Ethernet_LCD_HHPD), .PIN5(USB_HDMI_WiFi_BT_Ethernet_LCD_HHPD), .PIN4(USB_HDMI_WiFi_BT_Ethernet_LCD_HSDA), .PIN7(USB_HDMI_WiFi_BT_Ethernet_LCD_HSDA), .PIN10(USB_HDMI_WiFi_BT_Ethernet_LCD_HCEC), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_HCEC), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_HSCL), .PIN9(USB_HDMI_WiFi_BT_Ethernet_LCD_HSCL) );
  CELL_4_7k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R51 ( .PIN2(Net__HDMI1_Pad19_), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_HHPD) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R52 ( .PIN2(GND), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_HHPD) );
  BSS138_SOT23_3__OLIMEX_Transistors_FP_SOT23 FET1 ( .PIN1(_3_3VD), .PIN3(Net__FET1_Pad3_), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_HCEC) );
  CELL_27k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R46 ( .PIN1(_3_3VD), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_HCEC) );
  CELL_2_2k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R50 ( .PIN1(_5V), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_HSDA) );
  CELL_2_2k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R47 ( .PIN1(_5V), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_HSCL) );
  NA_510R__OLIMEX_RLC_FP_R_0402_5MIL_DWS R39 ( .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2P), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX2N) );
  NA_510R__OLIMEX_RLC_FP_R_0402_5MIL_DWS R43 ( .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1P), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX1N) );
  NA_510R__OLIMEX_RLC_FP_R_0402_5MIL_DWS R44 ( .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0P), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_HTX0N) );
  NA_510R__OLIMEX_RLC_FP_R_0402_5MIL_DWS R45 ( .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCP), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_HTXCN) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C79 ( .PIN1(GND), .PIN2(_3_3VD) );
  MICRO_USB_MISB_SWMM_5B_LF_OLIMEX_Connectors_FP_USB_MICRO_MISB_SWMM_5B_LF_Past USB_OTG1 ( .PIN0(GND), .PIN0(GND), .PIN0(GND), .PIN5(GND), .PIN0(GND), .PIN1(_5V_USBOTG), .PIN3(USB0_D_P), .PIN2(USB0_D_N), .PIN4(USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_ID) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R37 ( .PIN2(_3_3V), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_ID) );
  SY6280AAC_SOT23_5__OLIMEX_IC_FP_SOT_23_5 U6 ( .PIN2(GND), .PIN5(_5V), .PIN1(Net__C68_Pad2_), .PIN3(Net__R41_Pad2_), .PIN4(USB0_DRV) );
  FB0805_600R_2A_OLIMEX_RLC_FP_L_0805_5MIL_DWS L6 ( .PIN2(_5V_USBOTG), .PIN1(Net__C68_Pad2_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C67 ( .PIN2(GND), .PIN1(_5V_USBOTG) );
  NA_47uF_6_3V_20___OLIMEX_RLC_FP_C_0805_5MIL_DWS C70 ( .PIN1(GND), .PIN2(Net__C68_Pad2_) );
  NA_47uF_6_3V_20___OLIMEX_RLC_FP_C_0805_5MIL_DWS C69 ( .PIN1(GND), .PIN2(Net__C68_Pad2_) );
  CELL_47uF_6_3V_20__OLIMEX_RLC_FP_C_0805_5MIL_DWS C68 ( .PIN1(GND), .PIN2(Net__C68_Pad2_) );
  CELL_13k_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R41 ( .PIN1(GND), .PIN2(Net__R41_Pad2_) );
  CELL_4_7k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R38 ( .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_VBUSDET), .PIN2(Net__C68_Pad2_) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R42 ( .PIN1(GND), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_VBUSDET) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C72 ( .PIN1(GND), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_USB0_VBUSDET) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R40 ( .PIN1(GND), .PIN2(USB0_DRV) );
  CELL_47uF_6_3V_20__OLIMEX_RLC_FP_C_0805_5MIL_DWS C71 ( .PIN2(GND), .PIN1(_5V) );
  SY6280AAC_SOT23_5__OLIMEX_IC_FP_SOT_23_5 U9 ( .PIN2(GND), .PIN5(_5V), .PIN4(USB1_DRV), .PIN3(Net__R49_Pad2_), .PIN1(Net__C75_Pad2_) );
  FB0805_600R_2A_OLIMEX_RLC_FP_L_0805_5MIL_DWS L8 ( .PIN2(Net__C74_Pad1_), .PIN1(Net__C75_Pad2_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C74 ( .PIN2(GND), .PIN1(Net__C74_Pad1_) );
  NA_47uF_6_3V_20___OLIMEX_RLC_FP_C_0805_5MIL_DWS C77 ( .PIN1(GND), .PIN2(Net__C75_Pad2_) );
  NA_47uF_6_3V_20___OLIMEX_RLC_FP_C_0805_5MIL_DWS C76 ( .PIN1(GND), .PIN2(Net__C75_Pad2_) );
  CELL_47uF_6_3V_20__OLIMEX_RLC_FP_C_0805_5MIL_DWS C75 ( .PIN1(GND), .PIN2(Net__C75_Pad2_) );
  CELL_3_92k_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R49 ( .PIN1(GND), .PIN2(Net__R49_Pad2_) );
  NA_10k__OLIMEX_RLC_FP_R_0402_5MIL_DWS R48 ( .PIN1(GND), .PIN2(USB1_DRV) );
  CELL_47uF_6_3V_20__OLIMEX_RLC_FP_C_0805_5MIL_DWS C78 ( .PIN2(GND), .PIN1(_5V) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C73 ( .PIN1(GND), .PIN2(_3_3V) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C110 ( .PIN1(GND), .PIN2(_3_3VWiFiIO) );
  NA_RTL8723BS_ComboModule___OLIMEX_IC_FP_RL_SM02BD_RTL8723BS_ U11 ( .PIN31(GND), .PIN33(GND), .PIN36(GND), .PIN41(GND), .PIN1(GND), .PIN20(GND), .PIN9(_3_3V), .PIN22(_3_3VWiFiIO), .PIN34(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_RST_N), .PIN43(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_RX), .PIN38(Net__U11_Pad38_), .PIN29(Net__U11_Pad29_), .PIN3(Net__U11_Pad3_), .PIN30(Net__U11_Pad30_), .PIN32(Net__U11_Pad32_), .PIN35(Net__U11_Pad35_), .PIN37(Net__U11_Pad37_), .PIN23(Net__U11_Pad23_), .PIN39(Net__U11_Pad39_), .PIN4(Net__U11_Pad4_), .PIN40(Net__U11_Pad40_), .PIN5(Net__U11_Pad5_), .PIN6(USB_HDMI_WiFi_BT_Ethernet_LCD_AP_WAKE_BT), .PIN7(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_WAKE_AP), .PIN8(Net__U11_Pad8_), .PIN16(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_CMD), .PIN10(Net__U11_Pad10_), .PIN11(Net__U11_Pad11_), .PIN17(Net__R54_Pad1_), .PIN2(Net__C105_Pad1_), .PIN21(Net__U11_Pad21_), .PIN12(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_PMU_EN), .PIN13(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_WAKE_AP), .PIN42(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_TX), .PIN44(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_CTS), .PIN28(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_SYNC), .PIN26(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_CLK), .PIN27(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_DIN), .PIN25(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_PCM_DOUT), .PIN18(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D0), .PIN19(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D1), .PIN15(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D3), .PIN14(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D2), .PIN24(Net__R60_Pad1_) );
  NA_22R__OLIMEX_RLC_FP_R_0402_5MIL_DWS R54 ( .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_CLK), .PIN1(Net__R54_Pad1_) );
  NA_RA1206__4x0603__4B8_100k__OLIMEX_RLC_FP_RA1206__4X0603__4B8_xx RM9 ( .PIN4_1(_3_3VWiFiIO), .PIN3_1(_3_3VWiFiIO), .PIN2_1(_3_3VWiFiIO), .PIN1_1(_3_3VWiFiIO), .PIN4_2(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_PMU_EN), .PIN1_2(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D0), .PIN2_2(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D3), .PIN3_2(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D2) );
  NA_100nF_10V_10___OLIMEX_RLC_FP_C_0402_5MIL_DWS C92 ( .PIN1(GND), .PIN2(_3_3VWiFiIO) );
  NA_10uF_6_3V_20___OLIMEX_RLC_FP_C_0603_5MIL_DWS C91 ( .PIN1(GND), .PIN2(_3_3VWiFiIO) );
  NA_100nF_10V_10___OLIMEX_RLC_FP_C_0402_5MIL_DWS C90 ( .PIN1(GND), .PIN2(_3_3V) );
  NA_10uF_6_3V_20___OLIMEX_RLC_FP_C_0603_5MIL_DWS C89 ( .PIN1(GND), .PIN2(_3_3V) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C109 ( .PIN2(GND), .PIN1(VCC_PL) );
  NA_10pF_50V_5___OLIMEX_RLC_FP_C_0402_5MIL_DWS C105 ( .PIN1(Net__C105_Pad1_), .PIN2(Net__C105_Pad2_) );
  NA_0_8pF_C0402__OLIMEX_RLC_FP_C_0402_5MIL_DWS C106 ( .PIN1(GND), .PIN2(Net__C105_Pad2_) );
  NA_1_5pF_C0402__OLIMEX_RLC_FP_C_0402_5MIL_DWS C107 ( .PIN1(GND), .PIN2(Net__C107_Pad2_) );
  PCB_WIFI_ANT_OLIMEX_Antennas_FP_BT_Antenna_Inverted_1ANT_2GND ANT1 ( .PIN2(GND), .PIN1(Net__ANT1_Pad1_) );
  NA_RA1206__4x0603__4B8_100k__OLIMEX_RLC_FP_RA1206__4X0603__4B8_xx RM12 ( .PIN4_1(_3_3VWiFiIO), .PIN3_1(_3_3VWiFiIO), .PIN2_1(_3_3VWiFiIO), .PIN1_1(_3_3VWiFiIO), .PIN2_2(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_RST_N), .PIN4_2(USB_HDMI_WiFi_BT_Ethernet_LCD_BT_UART_RX), .PIN1_2(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_CMD), .PIN3_2(USB_HDMI_WiFi_BT_Ethernet_LCD_WL_SDIO_D1) );
  NA_10k__OLIMEX_RLC_FP_R_0402_5MIL_DWS R61 ( .PIN2(_3_3VWiFiIO), .PIN1(AP_CK32KO) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C80 ( .PIN2(GND), .PIN1(_3_3V) );
  CELL_2_2k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R70 ( .PIN2(_3_3V), .PIN1(TWI0_SCK) );
  CELL_2_2k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R71 ( .PIN2(_3_3V), .PIN1(TWI0_SDA) );
  FPV_WZA21_40_LF_OLIMEX_Connectors_FP_FPV_WZA21_40_LF LCD_CON1 ( .PIN22(GND), .PIN0(GND), .PIN13(GND), .PIN14(GND), .PIN2(GND), .PIN21(GND), .PIN4(GND), .PIN5(GND), .PIN6(GND), .PIN3(_3_3V), .PIN39(TWI0_SCK), .PIN40(TWI0_SDA), .PIN1(_5V), .PIN33(PH10), .PIN10(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD3_LCD_D21), .PIN20(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD0_LCD_D15), .PIN19(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD1_LCD_D14), .PIN18(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD2_LCD_D13), .PIN17(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD3_LCD_D12), .PIN8(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCTL_LCD_D19), .PIN31(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD0_LCD_CLK), .PIN11(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD2_LCD_D22), .PIN29(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCTL_LCD_HSYNC), .PIN36(USB_HDMI_WiFi_BT_Ethernet_LCD_GMDC_LCD_PWM), .PIN35(USB_HDMI_WiFi_BT_Ethernet_LCD_GMDIO_LCD_PWR), .PIN12(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD1_LCD_D23), .PIN9(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D20), .PIN15(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D10), .PIN16(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D11), .PIN23(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D2), .PIN24(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D3), .PIN25(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D4), .PIN26(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D5), .PIN27(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D6), .PIN28(USB_HDMI_WiFi_BT_Ethernet_LCD_LCD_D7), .PIN34(PH11), .PIN37(USB_HDMI_WiFi_BT_Ethernet_LCD_PH7_CTP_INT), .PIN32(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCK_LCD_DE), .PIN38(USB_HDMI_WiFi_BT_Ethernet_LCD_PH8_CTP_RST), .PIN30(USB_HDMI_WiFi_BT_Ethernet_LCD_GCLKIN_LCD_VSYNC), .PIN7(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCK_LCD_D18) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R99 ( .PIN1(_3_3V), .PIN2(USB1_DRV) );
  USB_A_VERTICAL_OLIMEX_Connectors_FP_USB_A_VERTICAL_PTH USB1 ( .PIN4(GND), .PIN0(GND), .PIN0(GND), .PIN1(Net__C74_Pad1_), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_USB1_DM), .PIN3(USB_HDMI_WiFi_BT_Ethernet_LCD_USB1_DP) );
  KSZ9031RNXCC_QFN48_1DRILL_PADPITCH_0_5MM___OLIMEX_IC_FP_QFN48_1DRILL_PADPITCH_0_5MM_ U15 ( .PIN49(GND), .PIN29(GND), .PIN48(Net__R115_Pad1_), .PIN33(Net__R105_Pad2_), .PIN41(Net__R109_Pad2_), .PIN47(Net__U15_Pad47_), .PIN38(Net__R119_Pad1_), .PIN43(Net__U15_Pad43_), .PIN46(Net__C212_Pad2_), .PIN10(USB_HDMI_WiFi_BT_Ethernet_LCD_MDI), .PIN15(Net__R113_Pad2_), .PIN12(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN34(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN40(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN16(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN13(Net__U15_Pad13_), .PIN17(Net__R111_Pad2_), .PIN45(Net__C213_Pad2_), .PIN42(Net__C211_Pad2_), .PIN22(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD3_LCD_D21), .PIN19(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD0_LCD_CLK), .PIN21(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD2_LCD_D22), .PIN25(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCTL_LCD_HSYNC), .PIN36(USB_HDMI_WiFi_BT_Ethernet_LCD_GMDC_LCD_PWM), .PIN37(USB_HDMI_WiFi_BT_Ethernet_LCD_GMDIO_LCD_PWR), .PIN20(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD1_LCD_D23), .PIN24(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCK_LCD_DE), .PIN35(Net__R107_Pad1_), .PIN44(Net__C207_Pad2_), .PIN4(Net__C207_Pad2_), .PIN9(Net__C207_Pad2_), .PIN14(Net__C204_Pad2_), .PIN39(Net__C204_Pad2_), .PIN30(Net__C204_Pad2_), .PIN18(Net__C204_Pad2_), .PIN23(Net__C204_Pad2_), .PIN26(Net__C204_Pad2_), .PIN28(Net__RM15_Pad3_1_), .PIN27(Net__RM15_Pad4_1_), .PIN31(Net__RM15_Pad2_1_), .PIN32(Net__RM15_Pad1_1_) );
  RA0805__4X0402__4_7k_OLIMEX_RLC_FP_RA0805__4X0402__xx_BIGGEROUTPADS RM8 ( .PIN1_1(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN2_1(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN4_1(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN3_1(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN3_2(Net__RM15_Pad3_1_), .PIN4_2(Net__RM15_Pad4_1_), .PIN2_2(Net__RM15_Pad2_1_), .PIN1_2(Net__RM15_Pad1_1_) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R105 ( .PIN2(Net__R105_Pad2_), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCTL_LCD_D19) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R106 ( .PIN2(Net__R105_Pad2_), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33) );
  CELL_1k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R107 ( .PIN2(GND), .PIN1(Net__R107_Pad1_) );
  NA_24pF_50V_5___OLIMEX_RLC_FP_C_0402_5MIL_DWS C198 ( .PIN2(Net__C198_Pad2_), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCK_LCD_D18) );
  CELL_1k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R108 ( .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_GMDIO_LCD_PWR) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R109 ( .PIN2(Net__R109_Pad2_), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_GCLKIN_LCD_VSYNC) );
  CELL_1k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R110 ( .PIN2(Net__R109_Pad2_), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33) );
  CELL_1k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R111 ( .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN2(Net__R111_Pad2_) );
  CELL_1k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R112 ( .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_PHYAD0), .PIN2(Net__R111_Pad2_) );
  CELL_1k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R113 ( .PIN2(Net__R113_Pad2_), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_PHYAD1) );
  CELL_1k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R114 ( .PIN1(GND), .PIN2(Net__R113_Pad2_) );
  TM211Q01FM22_OLIMEX_Connectors_FP_TM211Q01FM22 LAN1 ( .PIN9(USB_HDMI_WiFi_BT_Ethernet_LCD_MDI), .PIN14(USB_HDMI_WiFi_BT_Ethernet_LCD_PHYAD0), .PIN13(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN11(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN5(Net__C199_Pad2_), .PIN6(Net__C200_Pad2_), .SH2(Net__C196_Pad2_), .SH1(Net__C196_Pad2_), .PIN12(USB_HDMI_WiFi_BT_Ethernet_LCD_PHYAD1) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C199 ( .PIN1(GND), .PIN2(Net__C199_Pad2_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C200 ( .PIN1(GND), .PIN2(Net__C200_Pad2_) );
  CELL_1nF_2kV_10__X7R_OLIMEX_RLC_FP_C_1206_5MIL_DWS_ISO C196 ( .PIN1(GND), .PIN2(Net__C196_Pad2_) );
  FB0805_600R_2A_OLIMEX_RLC_FP_L_0805_5MIL_DWS L21 ( .PIN2(_3_3V), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33) );
  CELL_47uF_6_3V_20__OLIMEX_RLC_FP_C_0805_5MIL_DWS C201 ( .PIN2(GND), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C216 ( .PIN1(GND), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33) );
  CELL_22uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C214 ( .PIN1(GND), .PIN2(Net__C207_Pad2_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C207 ( .PIN1(GND), .PIN2(Net__C207_Pad2_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C215 ( .PIN1(GND), .PIN2(Net__C207_Pad2_) );
  CELL_47uF_6_3V_20__OLIMEX_RLC_FP_C_0805_5MIL_DWS C202 ( .PIN2(GND), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C217 ( .PIN1(GND), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C203 ( .PIN1(GND), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33) );
  CELL_22uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C204 ( .PIN1(GND), .PIN2(Net__C204_Pad2_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C208 ( .PIN1(GND), .PIN2(Net__C204_Pad2_) );
  CELL_22uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C205 ( .PIN1(GND), .PIN2(Net__C204_Pad2_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C209 ( .PIN1(GND), .PIN2(Net__C204_Pad2_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C206 ( .PIN1(GND), .PIN2(Net__C204_Pad2_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C210 ( .PIN1(GND), .PIN2(Net__C204_Pad2_) );
  CELL_12_1k_1__OLIMEX_RLC_FP_R_0603_5MIL_DWS R115 ( .PIN2(GND), .PIN1(Net__R115_Pad1_) );
  CELL_100k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R116 ( .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33), .PIN1(Net__C211_Pad2_) );
  CELL_1k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R117 ( .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_EPHY_RST_), .PIN1(Net__C211_Pad2_) );
  NA_OLIMEX_RLC_FP_R_0402_5MIL_DWS R118 ( .PIN2(AP_RESET_), .PIN1(Net__C211_Pad2_) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R119 ( .PIN1(Net__R119_Pad1_), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_VDD33) );
  CELL_1uF_10V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C211 ( .PIN1(GND), .PIN2(Net__C211_Pad2_) );
  CELL_27pF_50V_5__OLIMEX_RLC_FP_C_0402_5MIL_DWS C212 ( .PIN1(GND), .PIN2(Net__C212_Pad2_) );
  CELL_27pF_50V_5__OLIMEX_RLC_FP_C_0402_5MIL_DWS C213 ( .PIN1(GND), .PIN2(Net__C213_Pad2_) );
  FB0805_600R_2A_OLIMEX_RLC_FP_L_0805_5MIL_DWS L23 ( .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_1_25_EXT), .PIN1(Net__C207_Pad2_) );
  FB0805_600R_2A_OLIMEX_RLC_FP_L_0805_5MIL_DWS L24 ( .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_1_25_EXT), .PIN1(Net__C204_Pad2_) );
  CELL_22uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C218 ( .PIN2(GND), .PIN1(Net__C218_Pad1_) );
  AMS1117_ADJ__OLIMEX_Regulators_FP_SOT223 VR1 ( .PIN1(GND), .PIN3(Net__C218_Pad1_), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_1_25_EXT) );
  CELL_120R_OLIMEX_RLC_FP_R_0603_5MIL_DWS R120 ( .PIN2(GND), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_1_25_EXT) );
  CELL_22uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C219 ( .PIN2(GND), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_1_25_EXT) );
  HN1x2_Opened__OLIMEX_Jumpers_FP_HN1x2_Jumper PHYRST1 ( .PIN1(GND), .PIN2(Net__C211_Pad2_) );
  CELL_1N4007_SMA_OLIMEX_Diodes_FP_SMA_KA D5 ( .PIN2(_3_3V), .PIN1(Net__C218_Pad1_) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD CELL_1_25_EXT1 ( .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_1_25_EXT) );
  RA0805__4X0402__22R_OLIMEX_RLC_FP_RA0805__4X0402__xx_BIGGEROUTPADS RM15 ( .PIN1_2(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD0_LCD_D15), .PIN2_2(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD1_LCD_D14), .PIN3_2(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD2_LCD_D13), .PIN4_2(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXD3_LCD_D12), .PIN3_1(Net__RM15_Pad3_1_), .PIN4_1(Net__RM15_Pad4_1_), .PIN2_1(Net__RM15_Pad2_1_), .PIN1_1(Net__RM15_Pad1_1_) );
  RA0805__4X0402__22R_OLIMEX_RLC_FP_RA0805__4X0402__xx_BIGGEROUTPADS RM1 ( .PIN4_1(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD3_LCD_D21), .PIN2_1(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD0_LCD_CLK), .PIN3_1(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD2_LCD_D22), .PIN1_1(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXD1_LCD_D23), .PIN4_2(Net__RM1_Pad4_2_), .PIN1_2(Net__RM1_Pad1_2_), .PIN3_2(Net__RM1_Pad3_2_), .PIN2_2(Net__RM1_Pad2_2_) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R72 ( .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCTL_LCD_HSYNC), .PIN1(Net__R72_Pad1_) );
  NA_2_7nH_L0402__OLIMEX_RLC_FP_L_0402_5MIL_DWS L9 ( .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCK_LCD_DE), .PIN1(Net__C88_Pad2_) );
  NA_2_7nH_L0402__OLIMEX_RLC_FP_L_0402_5MIL_DWS L7 ( .PIN2(GND), .PIN1(Net__C198_Pad2_) );
  CELL_24pF_50V_5__OLIMEX_RLC_FP_C_0402_5MIL_DWS C93 ( .PIN1(GND), .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_GCLKIN_LCD_VSYNC) );
  NA_3_3nH___0_1nH_LQP15MN3N3B02D__OLIMEX_RLC_FP_L_0402_5MIL_DWS L10 ( .PIN2(Net__C105_Pad2_), .PIN1(Net__C107_Pad2_) );
  NA_24pF_50V_5___OLIMEX_RLC_FP_C_0402_5MIL_DWS C88 ( .PIN1(GND), .PIN2(Net__C88_Pad2_) );
  AT24C16C_SSHM_T_SOIC_8_150mil__OLIMEX_IC_FP_SOIC_8_150mil U4 ( .PIN4(GND), .PIN7(GND), .PIN2(_3_3V), .PIN3(_3_3V), .PIN8(_3_3V), .PIN1(_3_3V), .PIN5(TWI1_SDA), .PIN6(TWI1_SCK) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C39 ( .PIN2(GND), .PIN1(_3_3V) );
  NA_U_FL_R_SMT_1__OLIMEX_Connectors_FP_U_FL_R_SMT_1 ANT2 ( .PIN2(GND), .PIN1(Net__ANT2_Pad1_) );
  NA_0R__OLIMEX_RLC_FP_R_0402_5MIL_DWS R60 ( .PIN2(AP_CK32KO), .PIN1(Net__R60_Pad1_) );
  NA_0R__OLIMEX_RLC_FP_R_0402_5MIL_DWS R17 ( .PIN1(Net__ANT2_Pad1_), .PIN2(Net__C107_Pad2_) );
  CELL_0R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R16 ( .PIN2(Net__C107_Pad2_), .PIN1(Net__ANT1_Pad1_) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R18 ( .PIN2(Net__R107_Pad1_), .PIN1(USB_HDMI_WiFi_BT_Ethernet_LCD_GRXCK_LCD_D18) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R19 ( .PIN2(USB_HDMI_WiFi_BT_Ethernet_LCD_GTXCK_LCD_DE), .PIN1(Net__R19_Pad1_) );
  ABM8_25_000MHZ_D2Y_T_OLIMEX_Crystal_FP_TSX_3_2x2_5mm_GND_3_ Q4 ( .PIN3(GND), .PIN1(Net__C212_Pad2_), .PIN2(Net__C213_Pad2_) );
  CELL_1N5819_S4SOD_123__OLIMEX_Diodes_FP_SOD_123_1C_2A_KA D3 ( .PIN2(_5V), .PIN1(Net__D3_Pad1_) );
  ESDS314DBVR_SOT_23_5__OLIMEX_Diodes_FP_SOT_23_5 TVS1 ( .PIN2(GND) );
  ESDS314DBVR_SOT_23_5__OLIMEX_Diodes_FP_SOT_23_5 TVS2 ( .PIN2(GND), .PIN4(USB_HDMI_WiFi_BT_Ethernet_LCD_MDI) );
  AXP803_QFN68_8x8mm__OLIMEX_IC_FP_QFN68 U14 ( .PIN8(_1_5V), .PIN45(GND), .PIN69(GND), .PIN25(GND), .PIN12(GND), .PIN59(GND), .PIN20(_3_3V), .PIN68(_1_8V), .PIN31(_3_0VA), .PIN49(net_3_0V_RTC), .PIN28(VCC_PE), .PIN64(VBAT), .PIN46(AP_RESET_), .PIN1(Power_Supply__Extensions_and_MiPi_DSI_1_8V_DVDD_CSI), .PIN24(Net__U14_Pad24_), .PIN23(Net__U14_Pad23_), .PIN14(Power_Supply__Extensions_and_MiPi_DSI_2_8V_AVDD_CSI), .PIN16(Power_Supply__Extensions_and_MiPi_DSI_3_3V_MIPI), .PIN13(_3_3VWiFiIO), .PIN2(Net__C174_Pad2_), .PIN33(Net__C182_Pad2_), .PIN5(net_1_1V_CPUS), .PIN48(PMU_SDA), .PIN29(VCC_PL), .PIN27(Net__R87_Pad1_), .PIN26(Net__R86_Pad1_), .PIN65(Net__L18_Pad2_), .PIN34(Net__C151_Pad1_), .PIN35(Net__C149_Pad1_), .PIN30(Net__R83_Pad1_), .PIN53(Net__R82_Pad1_), .PIN41(VDDFB_CPUX), .PIN42(VDDFB_CPUX), .PIN62(Power_Supply__Extensions_and_MiPi_DSI_DC5SET), .PIN50(Net__C181_Pad2_), .PIN3(net_1_2V_HSIC), .PIN17(_3_3VD), .PIN9(net_1_1V_SYS), .PIN36(Net__L17_Pad1_), .PIN37(Net__L17_Pad1_), .PIN57(_5V_EXT), .PIN58(_5V_EXT), .PIN60(Net__C177_Pad2_), .PIN63(Net__C135_Pad1_), .PIN4(IPS), .PIN6(IPS), .PIN67(IPS), .PIN55(IPS), .PIN56(IPS), .PIN15(IPS), .PIN32(IPS), .PIN38(IPS), .PIN39(IPS), .PIN40(IPS), .PIN66(IPS), .PIN11(IPS), .PIN19(IPS), .PIN22(IPS), .PIN47(PMU_SCK), .PIN61(AP_NMI_), .PIN54(_5V_USBOTG), .PIN7(Net__L19_Pad1_), .PIN18(Net__C125_Pad2_), .PIN21(Net__L14_Pad1_), .PIN44(Net__L15_Pad1_), .PIN43(Net__L15_Pad1_), .PIN52(Net__T1_Pad3_), .PIN10(Net__L20_Pad1_), .PIN51(USB0_DRV) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C177 ( .PIN1(GND), .PIN2(Net__C177_Pad2_) );
  CELL_1k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R91 ( .PIN1(Net__PWRON1_Pad1_), .PIN2(Net__C177_Pad2_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C121 ( .PIN2(GND), .PIN1(_5V_EXT) );
  PWRJ_2mm_YDJ_1134__OLIMEX_Connectors_FP_PWRJ_2mm_YDJ_1134_ PWR1 ( ._(GND), ._(GND), ._(_5V_EXT) );
  NA_5025__OLIMEX_Devices_FP_FUSE_5025 FUSE2 ( .PIN1(_5V_EXT), .PIN2(_5V_EXT) );
  CELL_47uF_6_3V_20__OLIMEX_RLC_FP_C_0805_5MIL_DWS C118 ( .PIN1(GND), .PIN2(_5V_EXT) );
  CELL_47uF_6_3V_20__OLIMEX_RLC_FP_C_0805_5MIL_DWS C119 ( .PIN1(GND), .PIN2(_5V_EXT) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C124 ( .PIN2(GND), .PIN1(_5V_USBOTG) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C128 ( .PIN2(GND), .PIN1(IPS) );
  SWPA3015S1R5NT_1_5uH_2_30A_DCR_0_1R_CD32__OLIMEX_RLC_FP_CD32 L14 ( .PIN2(_3_3V), .PIN1(Net__L14_Pad1_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C122 ( .PIN1(GND), .PIN2(_3_3V) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C125 ( .PIN1(GND), .PIN2(Net__C125_Pad2_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C126 ( .PIN1(GND), .PIN2(IPS) );
  SWPA4018S1R5NT_1_5uH_3_35A_DCR_0_1R_CD43__OLIMEX_RLC_FP_CD42_43_ L15 ( .PIN2(net_1_1V_CPUX), .PIN1(Net__L15_Pad1_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C129 ( .PIN1(GND), .PIN2(net_1_1V_CPUX) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C131 ( .PIN1(GND), .PIN2(net_1_1V_CPUX) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C133 ( .PIN1(GND), .PIN2(IPS) );
  SWPA4018S1R5NT_1_5uH_3_35A_DCR_0_1R_CD43__OLIMEX_RLC_FP_CD42_43_ L17 ( .PIN1(Net__L17_Pad1_), .PIN2(net_1_1V_CPUX) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C136 ( .PIN1(GND), .PIN2(net_1_1V_CPUX) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C139 ( .PIN1(GND), .PIN2(net_1_1V_CPUX) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C145 ( .PIN1(GND), .PIN2(IPS) );
  SWPA3015S1R5NT_1_5uH_2_30A_DCR_0_1R_CD32__OLIMEX_RLC_FP_CD32 L19 ( .PIN2(_1_5V), .PIN1(Net__L19_Pad1_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C150 ( .PIN2(_1_5V), .PIN1(GND) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C153 ( .PIN1(GND), .PIN2(IPS) );
  NA_OLIMEX_RLC_FP_R_0402_5MIL_DWS R84 ( .PIN1(GND), .PIN2(Power_Supply__Extensions_and_MiPi_DSI_DC5SET) );
  SWPA3015S1R5NT_1_5uH_2_30A_DCR_0_1R_CD32__OLIMEX_RLC_FP_CD32 L20 ( .PIN2(net_1_1V_SYS), .PIN1(Net__L20_Pad1_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C154 ( .PIN1(GND), .PIN2(net_1_1V_SYS) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C157 ( .PIN1(GND), .PIN2(IPS) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C159 ( .PIN1(GND), .PIN2(IPS) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C161 ( .PIN1(GND), .PIN2(_3_3VD) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C162 ( .PIN1(GND), .PIN2(Power_Supply__Extensions_and_MiPi_DSI_3_3V_MIPI) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C164 ( .PIN1(GND), .PIN2(Power_Supply__Extensions_and_MiPi_DSI_2_8V_AVDD_CSI) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C165 ( .PIN1(GND), .PIN2(_3_3VWiFiIO) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C167 ( .PIN1(GND), .PIN2(IPS) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C176 ( .PIN1(GND), .PIN2(IPS) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C169 ( .PIN2(GND), .PIN1(IPS) );
  WPM1481_6_TR_DFN2X2_6L__OLIMEX_Transistors_FP_DFN2x2_6L T1 ( .PIN5(Net__C135_Pad1_), .PIN1(Net__C135_Pad1_), .PIN2(Net__C135_Pad1_), .PIN7(Net__C135_Pad1_), .PIN6(Net__C135_Pad1_), .PIN8(IPS), .PIN4(IPS), .PIN3(Net__T1_Pad3_) );
  CELL_0_01R_1__1206_OLIMEX_RLC_FP_R_1206_5MIL_DWS R78 ( .PIN2(VBAT), .PIN1(Net__C135_Pad1_) );
  CELL_1uF_10V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C135 ( .PIN2(VBAT), .PIN1(Net__C135_Pad1_) );
  SWPA4018S1R5NT_1_5uH_3_35A_DCR_0_1R_CD43__OLIMEX_RLC_FP_CD42_43_ L18 ( .PIN2(Net__L18_Pad2_), .PIN1(Net__C135_Pad1_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C144 ( .PIN2(GND), .PIN1(Net__C135_Pad1_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C138 ( .PIN2(GND), .PIN1(Net__C135_Pad1_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C147 ( .PIN2(GND), .PIN1(IPS) );
  LED_YELLOW_0603_OLIMEX_LEDs_FP_LED_0603_KA CHGLED1 ( .PIN1(Net__CHGLED1_Pad1_), .PIN2(IPS) );
  CELL_2_2k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R82 ( .PIN1(Net__R82_Pad1_), .PIN2(Net__CHGLED1_Pad1_) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R83 ( .PIN2(GND), .PIN1(Net__R83_Pad1_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C149 ( .PIN2(GND), .PIN1(Net__C149_Pad1_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C151 ( .PIN2(GND), .PIN1(Net__C151_Pad1_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C152 ( .PIN2(GND), .PIN1(net_3_0V_RTC) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R85 ( .PIN2(net_3_0V_RTC), .PIN1(AP_NMI_) );
  CELL_0R_Board_Mounted__OLIMEX_RLC_FP_R_0402_5MIL_0R_Board_Mounted_ R86 ( .PIN1(Net__R86_Pad1_), .PIN2(USB0_D_P) );
  CELL_0R_Board_Mounted__OLIMEX_RLC_FP_R_0402_5MIL_0R_Board_Mounted_ R87 ( .PIN1(Net__R87_Pad1_), .PIN2(USB0_D_N) );
  CELL_2_2k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R88 ( .PIN2(VCC_PL), .PIN1(PMU_SCK) );
  CELL_2_2k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R90 ( .PIN1(PMU_SDA), .PIN2(VCC_PL) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C173 ( .PIN2(GND), .PIN1(VCC_PL) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C175 ( .PIN2(GND), .PIN1(_3_0VA) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C171 ( .PIN2(GND), .PIN1(VCC_PE) );
  IT_1185AU2_160G_G_TR_OLIMEX_Buttons_FP_IT1185AU2_V2 PWRON1 ( .PIN2(GND), .PIN1(Net__PWRON1_Pad1_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C156 ( .PIN1(GND), .PIN2(AP_RESET_) );
  CELL_1k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R89 ( .PIN2(AP_RESET_), .PIN1(Net__R89_Pad1_) );
  IT_1185AU2_160G_G_TR_OLIMEX_Buttons_FP_IT1185AU2_V2 RESET1 ( .PIN2(GND), .PIN1(Net__R89_Pad1_) );
  CELL_1uF_10V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C160 ( .PIN1(GND), .PIN2(net_1_1V_SYS) );
  CELL_1uF_10V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C163 ( .PIN1(GND), .PIN2(net_1_1V_SYS) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C155 ( .PIN1(GND), .PIN2(net_1_1V_SYS) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C158 ( .PIN1(GND), .PIN2(net_1_1V_SYS) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C166 ( .PIN1(GND), .PIN2(net_1_1V_SYS) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C168 ( .PIN1(GND), .PIN2(net_1_1V_SYS) );
  CELL_1uF_10V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C142 ( .PIN1(GND), .PIN2(net_1_1V_CPUX) );
  CELL_1uF_10V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C137 ( .PIN1(GND), .PIN2(net_1_1V_CPUX) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C123 ( .PIN1(GND), .PIN2(net_1_1V_CPUX) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C148 ( .PIN1(GND), .PIN2(net_1_1V_CPUX) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C146 ( .PIN1(GND), .PIN2(net_1_1V_CPUX) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C127 ( .PIN1(GND), .PIN2(net_1_1V_CPUX) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C130 ( .PIN1(GND), .PIN2(net_1_1V_CPUX) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C132 ( .PIN1(GND), .PIN2(net_1_1V_CPUX) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C134 ( .PIN1(GND), .PIN2(net_1_1V_CPUX) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C117 ( .PIN1(GND), .PIN2(net_1_1V_CPUS) );
  CELL_1uF_10V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C120 ( .PIN1(GND), .PIN2(net_1_1V_CPUS) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C179 ( .PIN1(GND), .PIN2(net_1_1V_CPUS) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C115 ( .PIN1(GND), .PIN2(_3_3V) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C116 ( .PIN1(GND), .PIN2(_3_3V) );
  CELL_27pF_50V_5__OLIMEX_RLC_FP_C_0402_5MIL_DWS C185 ( .PIN2(GND), .PIN1(Net__C185_Pad1_) );
  CELL_27pF_50V_5__OLIMEX_RLC_FP_C_0402_5MIL_DWS C187 ( .PIN2(GND), .PIN1(Net__C187_Pad1_) );
  CELL_0R_Board_Mounted__OLIMEX_RLC_FP_R_0402_5MIL_0R_Board_Mounted_ R94 ( .PIN1(Net__R94_Pad1_), .PIN2(Net__C185_Pad1_) );
  Q32_768kHz_12_5pF_2P_SMD1206_OLIMEX_Crystal_FP_CM7V_T1A_Crystal_Package_1206_3_20x1_50x0_65mm_ Q2 ( .PIN1(Net__C183_Pad1_), .PIN2(Net__C184_Pad1_) );
  CELL_22pF_50V_5__OLIMEX_RLC_FP_C_0402_5MIL_DWS C183 ( .PIN2(GND), .PIN1(Net__C183_Pad1_) );
  CELL_22pF_50V_5__OLIMEX_RLC_FP_C_0402_5MIL_DWS C184 ( .PIN2(GND), .PIN1(Net__C184_Pad1_) );
  CELL_10M_OLIMEX_RLC_FP_R_0402_5MIL_DWS R93 ( .PIN1(Net__C183_Pad1_), .PIN2(Net__C184_Pad1_) );
  NA_OLIMEX_RLC_FP_R_0402_5MIL_DWS R96 ( .PIN2(GND), .PIN1(Net__R96_Pad1_) );
  NA_OLIMEX_RLC_FP_R_0402_5MIL_DWS R97 ( .PIN2(GND), .PIN1(Net__R97_Pad1_) );
  NA_OLIMEX_RLC_FP_R_0402_5MIL_DWS R98 ( .PIN2(GND), .PIN1(Net__R98_Pad1_) );
  NA_1nF_50V_10___OLIMEX_RLC_FP_C_0402_5MIL_DWS C193 ( .PIN1(GND), .PIN2(KEYADC) );
  IT_1185AU2_160G_G_TR_OLIMEX_Buttons_FP_IT1185AU2_V2 UBOOT1 ( .PIN2(GND), .PIN1(UBOOT) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C178 ( .PIN1(GND), .PIN2(net_1_2V_HSIC) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C186 ( .PIN1(GND), .PIN2(_3_3V) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C188 ( .PIN1(GND), .PIN2(Net__C188_Pad2_) );
  CELL_1uF_10V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C190 ( .PIN1(GND), .PIN2(net_3_0V_RTC) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C189 ( .PIN1(GND), .PIN2(net_3_0V_RTC) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C191 ( .PIN1(GND), .PIN2(_3_0VA) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C192 ( .PIN1(GND), .PIN2(Net__C192_Pad2_) );
  HN1x3_OLIMEX_Connectors_FP_HN1x3 DBG_UART1 ( .PIN3(GND), .PIN1(Net__DBG_UART1_Pad1_), .PIN2(Net__D4_Pad1_) );
  CELL_1N5819_S4SOD_123__OLIMEX_Diodes_FP_SOD_123_1C_2A_KA D4 ( .PIN1(Net__D4_Pad1_), .PIN2(Net__D4_Pad2_) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R95 ( .PIN2(_3_3V), .PIN1(Net__D4_Pad2_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C170 ( .PIN1(GND), .PIN2(_1_8V) );
  HN2x5_OLIMEX_Connectors_FP_HN2x5 UEXT1 ( .PIN2(GND), .PIN1(_3_3V), .PIN10(Power_Supply__Extensions_and_MiPi_DSI_UEXT_CS), .PIN3(UART3_TX), .PIN4(UART3_RX), .PIN6(TWI1_SDA), .PIN5(TWI1_SCK), .PIN8(Power_Supply__Extensions_and_MiPi_DSI_UEXT_MOSI), .PIN9(Power_Supply__Extensions_and_MiPi_DSI_UEXT_CLK), .PIN7(Power_Supply__Extensions_and_MiPi_DSI_UEXT_MISO) );
  CELL_2_2k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R75 ( .PIN1(_3_3V), .PIN2(TWI1_SCK) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R76 ( .PIN1(_3_3V), .PIN2(UART3_RX) );
  CELL_2_2k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R77 ( .PIN1(_3_3V), .PIN2(TWI1_SDA) );
  SMBJ6_0A_OLIMEX_Diodes_FP_DO214AA_1_K__2_A_ D1 ( .PIN2(GND), .PIN1(_5V_EXT) );
  LED_Red_0603_OLIMEX_LEDs_FP_LED_0603_KA PWRLED1 ( .PIN1(GND), .PIN2(Net__PWRLED1_Pad2_) );
  CELL_2_2k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R74 ( .PIN2(Net__PWRLED1_Pad2_), .PIN1(_5V_EXT) );
  Opened_OLIMEX_Jumpers_FP_SJ_1_SMALLER CELL_5V_E1 ( .PIN1(_5V_EXT), .PIN2(_5V) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C172 ( .PIN1(GND), .PIN2(Power_Supply__Extensions_and_MiPi_DSI_1_8V_DVDD_CSI) );
  NA_10uF_6_3V_20___OLIMEX_RLC_FP_C_0603_5MIL_DWS C174 ( .PIN1(GND), .PIN2(Net__C174_Pad2_) );
  CELL_1uF_10V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C181 ( .PIN1(GND), .PIN2(Net__C181_Pad2_) );
  CELL_1uF_10V_10__OLIMEX_RLC_FP_C_0603_5MIL_DWS C182 ( .PIN1(GND), .PIN2(Net__C182_Pad2_) );
  CELL_1k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R92 ( .PIN1(Power_Supply__Extensions_and_MiPi_DSI_DC5SET), .PIN2(Net__C181_Pad2_) );
  DW02R_OLIMEX_Connectors_FP_LIPO_BAT_CON2DW02R LIPO_BAT1 ( .PIN2(GND), .PIN1(VBAT) );
  CELL_47uF_6_3V_20__OLIMEX_RLC_FP_C_0805_5MIL_DWS C180 ( .PIN1(GND), .PIN2(VBAT) );
  NA_HN2x20__OLIMEX_Connectors_FP_HN2x20 GPIO1 ( .PIN2(GND), .PIN3(_3_3V), .PIN20(PC4), .PIN22(PC7), .PIN40(VCC_PE), .PIN34(PL12), .PIN24(PL7), .PIN26(PL8), .PIN28(PL9), .PIN30(PL10), .PIN32(PL11), .PIN6(UBOOT), .PIN31(Power_Supply__Extensions_and_MiPi_DSI_PE13), .PIN11(Power_Supply__Extensions_and_MiPi_DSI_PE3), .PIN9(Power_Supply__Extensions_and_MiPi_DSI_PE2), .PIN7(Power_Supply__Extensions_and_MiPi_DSI_PE1), .PIN5(Power_Supply__Extensions_and_MiPi_DSI_PE0), .PIN39(Power_Supply__Extensions_and_MiPi_DSI_PE17_GPIO_LED), .PIN35(Power_Supply__Extensions_and_MiPi_DSI_PE15), .PIN33(Power_Supply__Extensions_and_MiPi_DSI_PE14), .PIN13(Power_Supply__Extensions_and_MiPi_DSI_PE4), .PIN29(Power_Supply__Extensions_and_MiPi_DSI_PE12), .PIN27(Power_Supply__Extensions_and_MiPi_DSI_PE11), .PIN25(Power_Supply__Extensions_and_MiPi_DSI_PE10), .PIN23(Power_Supply__Extensions_and_MiPi_DSI_PE9), .PIN21(Power_Supply__Extensions_and_MiPi_DSI_PE8), .PIN19(Power_Supply__Extensions_and_MiPi_DSI_PE7), .PIN17(Power_Supply__Extensions_and_MiPi_DSI_PE6), .PIN15(Power_Supply__Extensions_and_MiPi_DSI_PE5), .PIN16(Power_Supply__Extensions_and_MiPi_DSI_PB3), .PIN14(Power_Supply__Extensions_and_MiPi_DSI_PB2), .PIN12(Power_Supply__Extensions_and_MiPi_DSI_PB1), .PIN10(Power_Supply__Extensions_and_MiPi_DSI_PB0), .PIN4(AP_RESET_), .PIN18(Power_Supply__Extensions_and_MiPi_DSI_PB4), .PIN36(Power_Supply__Extensions_and_MiPi_DSI_1_8V_DVDD_CSI), .PIN8(KEYADC), .PIN38(Power_Supply__Extensions_and_MiPi_DSI_2_8V_AVDD_CSI), .PIN1(_5V), .PIN37(Power_Supply__Extensions_and_MiPi_DSI_PE16_POWERON) );
  FPV_WZA21_20_LF_OLIMEX_Connectors_FP_FPV_WZA21_20_LF MIPI_DSI1 ( .PIN10(GND), .PIN1(GND), .PIN7(GND), .PIN18(GND), .PIN13(GND), .PIN4(GND), .PIN8(Power_Supply__Extensions_and_MiPi_DSI_DSI_D0N), .PIN15(Power_Supply__Extensions_and_MiPi_DSI_3_3V_MIPI), .PIN14(Power_Supply__Extensions_and_MiPi_DSI_3_3V_MIPI), .PIN11(TWI0_SCK), .PIN6(Power_Supply__Extensions_and_MiPi_DSI_DSI_CKP), .PIN16(Net__MIPI_DSI1_Pad16_), .PIN2(Power_Supply__Extensions_and_MiPi_DSI_DSI_D1N), .PIN3(Power_Supply__Extensions_and_MiPi_DSI_DSI_D1P), .PIN9(Power_Supply__Extensions_and_MiPi_DSI_DSI_D0P), .PIN5(Power_Supply__Extensions_and_MiPi_DSI_DSI_CKN), .PIN12(TWI0_SDA), .PIN19(Net__MIPI_DSI1_Pad19_), .PIN20(Net__MIPI_DSI1_Pad20_), .PIN17(Net__MIPI_DSI1_Pad17_) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C195 ( .PIN1(GND), .PIN2(_3_3V) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C194 ( .PIN1(GND), .PIN2(Net__3_3V_VCC_PE_2_8V1_Pad2_) );
  Opened_2_3__Closed_1_2__OLIMEX_Jumpers_FP_SJ_2_SMALL_12_TIED CELL_3_3V_VCC_PE_2_8V1 ( .PIN3(_3_3V), .PIN1(VCC_PE), .PIN2(Net__3_3V_VCC_PE_2_8V1_Pad2_) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R79 ( .PIN1(_3_3V), .PIN2(Power_Supply__Extensions_and_MiPi_DSI_UEXT_CS) );
  NA_2_2k__OLIMEX_RLC_FP_R_0402_5MIL_DWS R102 ( .PIN1(Power_Supply__Extensions_and_MiPi_DSI_PE15), .PIN2(Net__3_3V_VCC_PE_2_8V1_Pad2_) );
  NA_2_2k__OLIMEX_RLC_FP_R_0402_5MIL_DWS R101 ( .PIN1(Power_Supply__Extensions_and_MiPi_DSI_PE14), .PIN2(Net__3_3V_VCC_PE_2_8V1_Pad2_) );
  NA_B4B_PH_K_S__OLIMEX_Connectors_FP_B4B_PH_K_S HSIC1 ( .PIN4(GND), .PIN2(Net__HSIC1_Pad2_), .PIN3(Net__HSIC1_Pad3_), .PIN1(Net__HSIC1_Pad1_) );
  Opened_OLIMEX_Jumpers_FP_SJ HSIC_E1 ( .PIN2(Net__HSIC1_Pad1_), .PIN1(net_1_2V_HSIC) );
  CELL_100nF_10V_10__OLIMEX_RLC_FP_C_0402_5MIL_DWS C197 ( .PIN2(GND), .PIN1(net_1_2V_HSIC) );
  CELL_100k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R103 ( .PIN1(_3_0VA), .PIN2(KEYADC) );
  NA_10k__OLIMEX_RLC_FP_R_0402_5MIL_DWS R104 ( .PIN1(net_3_0V_RTC), .PIN2(AP_RESET_) );
  LED_Red_0603_OLIMEX_LEDs_FP_LED_0603_KA GPIO_LED1 ( .PIN1(GND), .PIN2(Net__GPIO_LED1_Pad2_) );
  CELL_1k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R58 ( .PIN2(Net__GPIO_LED1_Pad2_), .PIN1(Power_Supply__Extensions_and_MiPi_DSI_PE17_GPIO_LED) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD CELL_3_3V1 ( .PIN1(_3_3V) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD CELL_1_1V_CPUX1 ( .PIN1(net_1_1V_CPUX) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD DDR_VCC1 ( .PIN1(_1_5V) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD CELL_1_1V_SYS1 ( .PIN1(net_1_1V_SYS) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD _3_3VD1 ( .PIN1(_3_3VD) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD _3_3VWiFiIO1 ( .PIN1(_3_3VWiFiIO) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD CELL_3_3V_MIPI1 ( .PIN1(Power_Supply__Extensions_and_MiPi_DSI_3_3V_MIPI) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD _5V_USBOTG1 ( .PIN1(_5V_USBOTG) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD IPS1 ( .PIN1(IPS) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD CELL_3_0V_RTC1 ( .PIN1(net_3_0V_RTC) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD VCC_PC1 ( .PIN1(VCC_PC) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD _1_8V1 ( .PIN1(_1_8V) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD CELL_1_1V_CPUS1 ( .PIN1(net_1_1V_CPUS) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD _3_0VA1 ( .PIN1(_3_0VA) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD VCC_PL1 ( .PIN1(VCC_PL) );
  TESTPAD_OLIMEX_TestPoints_FP_TP_SMD GND1 ( .PIN1(GND) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R65 ( .PIN2(Power_Supply__Extensions_and_MiPi_DSI_PE16), .PIN1(Power_Supply__Extensions_and_MiPi_DSI_PE16_POWERON) );
  NA_1k__OLIMEX_RLC_FP_R_0402_5MIL_DWS R28 ( .PIN2(Net__C177_Pad2_), .PIN1(Power_Supply__Extensions_and_MiPi_DSI_PE16_POWERON) );
  Opened_2_3__Soldered_1_2__OLIMEX_Jumpers_FP_SJ_2_SMALL PWR_PC1 ( .PIN1(_3_3V), .PIN3(_1_8V), .PIN2(VCC_PC) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R121 ( .PIN2(SPI0_MISO), .PIN1(Power_Supply__Extensions_and_MiPi_DSI_UEXT_MISO) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R122 ( .PIN2(SPI0_CLK), .PIN1(Power_Supply__Extensions_and_MiPi_DSI_UEXT_CLK) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R123 ( .PIN1(SPI0_MOSI), .PIN2(Power_Supply__Extensions_and_MiPi_DSI_UEXT_MOSI) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R124 ( .PIN1(SPI0_CS), .PIN2(Power_Supply__Extensions_and_MiPi_DSI_UEXT_CS) );
  NA_22R__OLIMEX_RLC_FP_R_0402_5MIL_DWS R73 ( .PIN2(Power_Supply__Extensions_and_MiPi_DSI_UEXT_CS), .PIN1(PH10) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R125 ( .PIN2(Power_Supply__Extensions_and_MiPi_DSI_DSI_D3P), .PIN1(Net__MIPI_DSI1_Pad17_) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R126 ( .PIN2(Power_Supply__Extensions_and_MiPi_DSI_DSI_D2N), .PIN1(Net__MIPI_DSI1_Pad19_) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R130 ( .PIN1(Power_Supply__Extensions_and_MiPi_DSI_DSI_D2P), .PIN2(Net__MIPI_DSI1_Pad20_) );
  CELL_22R_OLIMEX_RLC_FP_R_0402_5MIL_DWS R129 ( .PIN1(Power_Supply__Extensions_and_MiPi_DSI_DSI_D3N), .PIN2(Net__MIPI_DSI1_Pad16_) );
  NA_OLIMEX_RLC_FP_R_0402_5MIL_DWS R128 ( .PIN2(Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_EN), .PIN1(Net__MIPI_DSI1_Pad19_) );
  NA_OLIMEX_RLC_FP_R_0402_5MIL_DWS R127 ( .PIN2(Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_RST), .PIN1(Net__MIPI_DSI1_Pad17_) );
  NA_OLIMEX_RLC_FP_R_0402_5MIL_DWS R132 ( .PIN1(Power_Supply__Extensions_and_MiPi_DSI_MIPI_DSI_BKL), .PIN2(Net__MIPI_DSI1_Pad20_) );
  NA_OLIMEX_RLC_FP_R_0402_5MIL_DWS R131 ( .PIN2(Net__MIPI_DSI1_Pad16_), .PIN1(IPS) );
  ABM8_24_000MHZ_D2Y_T_OLIMEX_Crystal_FP_TSX_3_2x2_5mm_GND_3_ Q3 ( .PIN3(GND), .PIN2(Net__C187_Pad1_), .PIN1(Net__C185_Pad1_) );
  VDA4510CTA_SOT_23__OLIMEX_IC_FP_SOT_23 U16 ( .PIN2(GND), .PIN3(_5V_EXT), .PIN1(Net__FET3_Pad1_) );
  BSS138_SOT23_3__OLIMEX_Transistors_FP_SOT23 FET4 ( .PIN2(GND), .PIN1(Net__FET3_Pad1_), .PIN3(Net__FET2_Pad1_) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R20 ( .PIN2(_5V_EXT), .PIN1(Net__FET3_Pad1_) );
  CELL_10k_OLIMEX_RLC_FP_R_0402_5MIL_DWS R24 ( .PIN2(Net__FET2_Pad1_), .PIN1(_5V) );
  IRLML6402_SOT_23__OLIMEX_Transistors_FP_SOT23 FET2 ( .PIN3(_5V_EXT), .PIN1(Net__FET2_Pad1_), .PIN2(_5V) );
  CELL_1M_OLIMEX_RLC_FP_R_0402_5MIL_DWS R22 ( .PIN1(GND), .PIN2(Net__FET3_Pad1_) );
  IRLML6402_SOT_23__OLIMEX_Transistors_FP_SOT23 FET3 ( .PIN1(Net__FET3_Pad1_), .PIN2(_5V), .PIN3(Net__C143_Pad2_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C143 ( .PIN1(GND), .PIN2(Net__C143_Pad2_) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C140 ( .PIN1(GND), .PIN2(IPS) );
  CELL_1_1k_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R81 ( .PIN2(GND), .PIN1(Net__R80_Pad2_) );
  CELL_8_25k_1__OLIMEX_RLC_FP_R_0402_5MIL_DWS R80 ( .PIN1(Net__C143_Pad2_), .PIN2(Net__R80_Pad2_) );
  CELL_1N5822_SS34_SMA_OLIMEX_Diodes_FP_SMA_KA D2 ( .PIN2(Net__D2_Pad2_), .PIN1(Net__C143_Pad2_) );
  CELL_2_2uH_3A_YS75_7x8_OLIMEX_RLC_FP_YS75_7X8MM L16 ( .PIN2(Net__D2_Pad2_), .PIN1(IPS) );
  CELL_10uF_6_3V_20__OLIMEX_RLC_FP_C_0603_5MIL_DWS C141 ( .PIN1(GND), .PIN2(IPS) );
  MT3608_SOT23_6__OLIMEX_IC_FP_SOT23_6 U13 ( .PIN2(GND), .PIN4(_3_3V), .PIN1(Net__D2_Pad2_), .PIN3(Net__R80_Pad2_), .PIN6(Net__U13_Pad6_), .PIN5(IPS) );
endmodule